// Build a circuit with no inputs and one output that outputs a constant 0

module top_module(
    output zero
);// Module body starts after semicolon

    assign zero = 0;
    
endmodule

